module RegFile (
    input  logic         clk,
    input  logic         rst,
    input  logic  [4:0]  rs1_addr,
    input  logic  [4:0]  rs2_addr,
    input  logic  [4:0]  rd_addr,
    input  logic  [31:0] rd_data,
    input  logic         rd_we,
    output logic [31:0]  rs1_data,
    output logic [31:0]  rs2_data
);

    logic [31:0] regs [31:0];

    // Read ports
    assign rs1_data = (rs1_addr == 0) ? 32'b0 : regs[rs1_addr];
    assign rs2_data = (rs2_addr == 0) ? 32'b0 : regs[rs2_addr];

    // Write port
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            regs <= '{default:32'b0};
        end else if (rd_we && (rd_addr != 0)) begin
            regs[rd_addr] <= rd_data;
        end
    end

endmodule